// ============================================================================
// Designer : Yi_Yuan Chen
// Create   : 2022.12.09
// Ver      : 1.0
// Func     : output top module
// 			Unsupport output channel less than 8.
// 			If change PE block number parameter !=8 , plz check all module connection 
// 			cause paramize is not ready.
// ============================================================================
//      Instance Name:              OT_SRAM
//      Words:                      1024
//      Bits:                       64
//      Mux:                        8
//      Drive:                      6
//      Write Mask:                 Off
//      Extra Margin Adjustment:    On
//      Accelerated Retention Test: Off
//      Redundant Rows:             0
//      Redundant Columns:          0
//      Test Muxes                  Off
//----------------------------------------------------------------------------------
//                   /--------------  output top  --------------------------------------------------------\
//	/----------\  -> | /---------------\  -> /-----------\     /---------\     /----------\    /---------\|
//	| PEblk_n..| --> | | qtbuf_mod_n.. | --> |  bit_mux  | --> | qtbfifo | --> | ot_write | -->| ot_read ||   
//	\----------/  -> | \---------------/  -> \-----------/     \---------/     \----------/    \---------/|
//                   \--------------  output top  --------------------------------------------------------/
//--------------------------------------------------------------------------------


module ot_top 
#(
	parameter TBITS = 64 
	,	TBYTE = 8
	,	PEBLKROW_NUM = 8
	,	SRAM_DATA_BITS = 64
	,	SRAM_ADDR_BITS = 10
)(
	clk 	
	,	reset 				

	,	fifo_full_n			
	,	fifo_write			
	,	fifo_last			
	,	fifo_data			

	,	valid_din 			
	,	data_din		

	,	cfg_ot_rnd_finsub1	
	,	cfg_ot_tgpfnsub1	
	,	cfg_ot_tcolfnsub1	
	,	cfg_ot_tchafnsub1	
	,	cfg_ot_sft_gp		
	,	cfg_ot_sft_colpra	
);
	

	// localparam SRAM_DATA_BITS = 64;
	// localparam SRAM_ADDR_BITS = 10;

//==============================================================================
//========    I/O Signal Declare    ========
//==============================================================================

	input clk		;
	input reset		;

	input [ PEBLKROW_NUM-1:0]			valid_din		;
	input [ PEBLKROW_NUM*TBITS-1 : 0 ]		data_din		;

	input 	fifo_full_n		;
	output	fifo_write		;
	output	fifo_last		;
	output [ SRAM_DATA_BITS-1 : 0 ]	fifo_data		;
	
	//----    config in    -----
	input wire	[ SRAM_ADDR_BITS-1 : 0 ]	cfg_ot_rnd_finsub1	;
	input wire	[ SRAM_ADDR_BITS-1 : 0 ]	cfg_ot_tgpfnsub1	;
	input wire	[ SRAM_ADDR_BITS-1 : 0 ]	cfg_ot_tcolfnsub1	;
	input wire	[ SRAM_ADDR_BITS-1 : 0 ]	cfg_ot_tchafnsub1	;
	input wire	[ SRAM_ADDR_BITS-1 : 0 ]	cfg_ot_sft_gp		;
	input wire	[ SRAM_ADDR_BITS-1 : 0 ]	cfg_ot_sft_colpra	;
//-----------------------------------------------------------------------------

//==============================================================================
//========    output module config register    ========
//==============================================================================

reg [ SRAM_ADDR_BITS-1 : 0 ]	rcfg_ot_rnd_finsub1 ;
reg [ SRAM_ADDR_BITS-1 : 0 ]	rcfg_ot_tgpfnsub1	;
reg [ SRAM_ADDR_BITS-1 : 0 ]	rcfg_ot_tcolfnsub1	;
reg [ SRAM_ADDR_BITS-1 : 0 ]	rcfg_ot_tchafnsub1	;
reg [ SRAM_ADDR_BITS-1 : 0 ]	rcfg_ot_sft_gp		;
reg [ SRAM_ADDR_BITS-1 : 0 ]	rcfg_ot_sft_colpra	;

//-----------------------------------------------------------------------------
//----    temporal cfg setting    -----
always @(posedge clk ) begin
	if(reset)begin
		rcfg_ot_rnd_finsub1 <= 191	;
		rcfg_ot_tgpfnsub1	<= 1	;
		rcfg_ot_tcolfnsub1	<= 7	;
		rcfg_ot_tchafnsub1	<= 7	;
		rcfg_ot_sft_gp		<= 64	;
		rcfg_ot_sft_colpra	<= 8	;
	end
	else begin
		rcfg_ot_rnd_finsub1 <= cfg_ot_rnd_finsub1	;
		rcfg_ot_tgpfnsub1	<= cfg_ot_tgpfnsub1	;
		rcfg_ot_tcolfnsub1	<= cfg_ot_tcolfnsub1	;
		rcfg_ot_tchafnsub1	<= cfg_ot_tchafnsub1	;
		rcfg_ot_sft_gp		<= cfg_ot_sft_gp		;
		rcfg_ot_sft_colpra	<= cfg_ot_sft_colpra	;
	end
end
//-----------------------------------------------------------------------------
//-----------------------------------------------------------------------------


//----generated by ot_top_mod.py------ 
//---- ot_top declare OT_SRAM start------ 
wire cen_otsr_0 ,cen_otsr_1 ; 
wire wen_otsr_0 ,wen_otsr_1 ; 
wire [ SRAM_ADDR_BITS -1 : 0 ] addr_otsr_0 ,addr_otsr_1 ; 
wire [ SRAM_DATA_BITS -1 : 0 ] din_otsr_0 ,din_otsr_1 ; 
wire [ SRAM_DATA_BITS -1 : 0 ] dout_otsr_0 ,dout_otsr_1 ; 
//---- ot top declare OT_SRAM end------ 


//----declare ot_top sram read signal start------ 
wire osr_cen_otsr_0 ; 
wire osr_wen_otsr_0 ; 
wire [ SRAM_ADDR_BITS -1 : 0 ] osr_addr_otsr_0 ; 
wire [ SRAM_DATA_BITS -1 : 0 ] osr_dout_otsr_0 ; 
//----declare ot_top sram read signal  end------ 


//----declare ot_top sram write signal start------ 
wire osw_cen_otsr_0 ; 
wire osw_wen_otsr_0 ; 
wire [ SRAM_ADDR_BITS -1 : 0 ] osw_addr_otsr_0 ; 
wire [ SRAM_DATA_BITS -1 : 0 ] osw_din_otsr_0 ; 
//----declare ot_top sram write signal  end------ 


localparam BUF_STATE_BITS = 3;
localparam IDLE 	= 3'd0;
localparam READY 	= 3'd1;

localparam WRING 	= 3'd2;
localparam WR_DONE 	= 3'd3;
localparam RDING 	= 3'd4;
localparam RD_DONE 	= 3'd5;

reg [BUF_STATE_BITS-1: 0 ] bf0_current_state ;
reg [BUF_STATE_BITS-1: 0 ] bf0_next_state ;

reg [BUF_STATE_BITS-1: 0 ] bf1_current_state ;
reg [BUF_STATE_BITS-1: 0 ] bf1_next_state ;


wire write_last ;
wire dual_done ;

reg read_start ;
wire read_busy ;
wire read_done ;

//------- qtb and fifo signal --------
wire fifo_empty_n 	;
wire fifo_read 		;
wire valid_2_otfifo	;
wire [ TBITS-1 : 0 ]data64_2_otfifo	;
wire [ TBITS-1 : 0 ] fifo_data64	;
wire fifo_w_empty_n	;
wire fifo_w_read	;
//-----------------------------------------------------------------------------
//----    qtb Declare    -----
wire [TBITS-1:0]	qtb_qresult	[0:PEBLKROW_NUM-1]	;
wire			qtb_qvalid	[0:PEBLKROW_NUM-1]	;
wire [ TBITS-1 : 0 ]	qtb_64bitsout	[0:PEBLKROW_NUM-1]	;
wire			qtb_validout	[0:PEBLKROW_NUM-1]	;
//-----------------------------------------------------------------------------
//----    bit mux Declare    -----
wire [PEBLKROW_NUM-1:0]					qtb2bitmux_valid	;
wire [PEBLKROW_NUM*TBITS -1 : 0]		qtb2bitmux_data		;
//-----------------------------------------------------------------------------
//----    actually cen wen signal declare    -----
wire atl_cen_otsr_0 ;	// for actually connection between FPGA and CBDK
wire atl_wen_otsr_0 ;	// for actually connection between FPGA and CBDK
wire atl_cen_otsr_1 ;	// for actually connection between FPGA and CBDK
wire atl_wen_otsr_1 ;	// for actually connection between FPGA and CBDK
//-----------------------------------------------------------------------------

// =============================================================================
// ========================    SRAM instance     ===============================
// =============================================================================
`ifdef FPGA_SRAM_SETTING
	BRAM_OT otbf_0 ( .clka( clk ) ,.ena( atl_cen_otsr_0 )	,.wea( atl_wen_otsr_0 )	,.addra( addr_otsr_0 ),.dina( din_otsr_0 )	,.douta( dout_otsr_0 ) );
	BRAM_OT otbf_1 ( .clka( clk ) ,.ena( atl_cen_otsr_1 )	,.wea( atl_wen_otsr_1 )	,.addra( addr_otsr_1 ),.dina( din_otsr_1 )	,.douta( dout_otsr_1 ) );
`else 
	//----generated by ot_top_mod.py------ 
	//----instance OT_SRAM start------ 
	OT_SRAM otbf_0(.Q(	dout_otsr_0 ),	.CLK( clk ),.CEN( atl_cen_otsr_0 ),.WEN( atl_wen_otsr_0 ),.A( addr_otsr_0 ),.D( din_otsr_0 ),.EMA( 3'b0 ));//----instance OT SRAM_0---------
	OT_SRAM otbf_1(.Q(	dout_otsr_1 ),	.CLK( clk ),.CEN( atl_cen_otsr_1 ),.WEN( atl_wen_otsr_1 ),.A( addr_otsr_1 ),.D( din_otsr_1 ),.EMA( 3'b0 ));//----instance OT SRAM_1---------
	//----instance OT_SRAM end------ 
`endif 
// //----generated by ot_top_mod.py------ 
// //----instance OT_SRAM start------ 
// OT_SRAM otbf_0(.Q(	dout_otsr_0 ),	.CLK( clk ),.CEN( cen_otsr_0 ),.WEN( wen_otsr_0 ),.A( addr_otsr_0 ),.D( din_otsr_0 ),.EMA( 3'b0 ));//----instance OT SRAM_0---------
// OT_SRAM otbf_1(.Q(	dout_otsr_1 ),	.CLK( clk ),.CEN( cen_otsr_1 ),.WEN( wen_otsr_1 ),.A( addr_otsr_1 ),.D( din_otsr_1 ),.EMA( 3'b0 ));//----instance OT SRAM_1---------
// //----instance OT_SRAM end------ 


//-----------------------------------------------------------------------------


// ===============================================================
// ==============		ot module instance		==================
// ===============================================================
ot_write #(
	.SRAM_DATA_BITS( SRAM_DATA_BITS )
	,	.SRAM_ADDR_BITS( SRAM_ADDR_BITS )
)ow000 (
	.clk			(	clk				)
	,	.reset			(	reset			)
	,	.data_in		(	fifo_data64			)
	,	.fifo_empty_n	(	fifo_w_empty_n	)
	,	.fifo_read 		(	fifo_w_read	)

	,	.last			(	write_last		)
	,	.cen_otsr		(	osw_cen_otsr_0		)
	,	.wen_otsr		(	osw_wen_otsr_0		)
	,	.addr_otsr		(	osw_addr_otsr_0		)
	,	.data_for_sram	(	osw_din_otsr_0		)
	,	.cfg_ot_rnd_finsub1	(	rcfg_ot_rnd_finsub1		)

);

ot_read #(
	.SRAM_DATA_BITS( SRAM_DATA_BITS )
	,	.SRAM_ADDR_BITS( SRAM_ADDR_BITS )
)
or111 (
	.clk			(	clk				)
	,	.reset			(	reset			)

	,	.start			(	read_start	)
	,	.busy			(	read_busy	)
	,	.done			(	read_done	)
	,	.fifo_full_n	(	fifo_full_n	)
	,	.fifo_write		(	fifo_write	)
	,	.fifo_last		(	fifo_last	)
	,	.fifo_data		(	fifo_data	)

	,	.data_from_sram	(	osr_dout_otsr_0	)
	,	.addr_otsr		(	osr_addr_otsr_0	)
	,	.cen_otsr		(	osr_cen_otsr_0	)
	,	.wen_otsr		(	osr_wen_otsr_0	)


	,	.cfg_ot_tgpfnsub1	(	rcfg_ot_tgpfnsub1		)
	,	.cfg_ot_tcolfnsub1	(	rcfg_ot_tcolfnsub1		)
	,	.cfg_ot_tchafnsub1	(	rcfg_ot_tchafnsub1		)
	,	.cfg_ot_sft_gp		(	rcfg_ot_sft_gp			)
	,	.cfg_ot_sft_colpra	(	rcfg_ot_sft_colpra		)

);


ot_fifo  qtbfifo(
	.clk			(	clk		),
	.reset			(	reset	),
	.valid_in 		(	valid_2_otfifo	),
	.data_in		(	data64_2_otfifo	),
	// .error			(		),	// we loss output data cause something wrong
	.empty_n		(	fifo_empty_n	),
	.read			(	fifo_read		),
	.data_out		(	fifo_data64		)
);


ot_bitmux64 #(
	.TBITS (TBITS )
	,	.PEBLKROW_NUM  ( PEBLKROW_NUM )
)dd(
	.clk 			(	clk		)
	,	.reset 			(	reset	)
	,	.valid_din 		(	{ qtb_qvalid[0] , qtb_qvalid[1] , qtb_qvalid[2] , qtb_qvalid[3] , qtb_qvalid[4] , qtb_qvalid[5] , qtb_qvalid[6] , qtb_qvalid[7] }	)
	,	.data_din		(	{ qtb_qresult[0] , qtb_qresult[1] , qtb_qresult[2] , qtb_qresult[3] , qtb_qresult[4] , qtb_qresult[5] , qtb_qresult[6] , qtb_qresult[7] }		)
	,	.valid_dout		(	valid_2_otfifo	)
	,	.result_dout		(	data64_2_otfifo	)
);

//----    quan to buffer module instance    -----
// genvar gx ;
// generate
// 	for(gx=0; gx< PEBLKROW_NUM ; gx=gx+1)begin	: inst_qtb
// 		ot_qtbuf	qtb0(
// 			.clk				(	clk		)
// 			,	.reset 			(	reset		)
// 			,	.q_result_din	(	qtb_qresult[gx]		)
// 			,	.q_valid_din	(	qtb_qvalid[gx]		)
// 			,	.out64bits		(	qtb_64bitsout[gx]	)
// 			,	.valid_out		(	qtb_validout[gx]	)
// 		);
// 	end
// endgenerate
// ot_qtbuf	qtb00(
// 	.clk				(	clk		)
// 	,	.reset 			(	reset		)
// 	,	.q_result_din	(	qtb_qresult[gx]		)
// 	,	.q_valid_din	(	qtb_qvalid[gx]	)
	
// 	,	.out64bits		(	qtb_64bitsout[gx]	)
// 	,	.valid_out		(	qtb_validout[gx]	)

// );
//-----------------------------------------------------------------------------


assign qtb2bitmux_valid = {
		qtb_validout[0]
		,	qtb_validout[1]
		,	qtb_validout[2]
		,	qtb_validout[3]
		,	qtb_validout[4]
		,	qtb_validout[5]
		,	qtb_validout[6]
		,	qtb_validout[7]
};
assign qtb2bitmux_data = {
		qtb_64bitsout[0]
		,	qtb_64bitsout[1]
		,	qtb_64bitsout[2]
		,	qtb_64bitsout[3]
		,	qtb_64bitsout[4]
		,	qtb_64bitsout[5]
		,	qtb_64bitsout[6]
		,	qtb_64bitsout[7]
};





genvar gy ;
generate
	for (gy = 0; gy<PEBLKROW_NUM; gy=gy+1) begin	:assq_result
		assign	qtb_qresult[gy] = data_din[ (TBITS*(PEBLKROW_NUM-gy)-1)	-:	TBITS	] ;
		assign	qtb_qvalid[gy] = valid_din[ (PEBLKROW_NUM-1 -gy)	-:	1	] ;
	end
endgenerate



`ifdef FPGA_SRAM_SETTING
	assign atl_cen_otsr_0 	= ~cen_otsr_0;
	assign atl_wen_otsr_0 	= ~wen_otsr_0;
	assign atl_cen_otsr_1 	= ~cen_otsr_1;
	assign atl_wen_otsr_1 	= ~wen_otsr_1;
`else 
	assign atl_cen_otsr_0 	= cen_otsr_0	;
	assign atl_wen_otsr_0 	= wen_otsr_0	;
	assign atl_cen_otsr_1 	= cen_otsr_1	;
	assign atl_wen_otsr_1 	= wen_otsr_1	;
`endif 

assign cen_otsr_0 	= ( bf0_current_state == WRING )? osw_cen_otsr_0 : 
						( bf0_current_state == RDING )? osr_cen_otsr_0 : 1'd1 	;
assign wen_otsr_0 	= ( bf0_current_state == WRING )? osw_wen_otsr_0 :  1'd1 	;
assign din_otsr_0 	= osw_din_otsr_0	;
assign addr_otsr_0	= ( bf0_current_state == WRING )? osw_addr_otsr_0 : 
						( bf0_current_state == RDING )? osr_addr_otsr_0 : 10'd0 	;

assign cen_otsr_1 	= ( bf1_current_state == WRING )? osw_cen_otsr_0 : 
						( bf1_current_state == RDING )? osr_cen_otsr_0 : 1'd1 	;
assign wen_otsr_1 	= ( bf1_current_state == WRING )? osw_wen_otsr_0 :  1'd1 	;
assign din_otsr_1 	= osw_din_otsr_0	;
assign addr_otsr_1	= ( bf1_current_state == WRING )? osw_addr_otsr_0 : 
						( bf1_current_state == RDING )? osr_addr_otsr_0 : 10'd0 	;


assign osr_dout_otsr_0 = ( bf0_current_state == RDING )? dout_otsr_0 :
							( bf1_current_state == RDING )? dout_otsr_1 :	64'd0 ;




assign fifo_w_empty_n = (  (bf0_current_state == WRING ) | ( bf1_current_state == WRING ) ) ? fifo_empty_n : 1'd0 ;
assign fifo_read = (  (bf0_current_state == WRING ) | ( bf1_current_state == WRING ) ) ? 	fifo_w_read : 1'd0 ;






//==============================================================================
//========    Buffer read/write control    ========
//==============================================================================
always @(posedge clk ) begin
	if(reset )begin
		bf0_current_state <= WRING ;
		bf1_current_state <= IDLE ;
	end
	else begin
		bf0_current_state <= bf0_next_state ;
		bf1_current_state <= bf1_next_state ;
	end
end


always @(*) begin
	case (bf0_current_state)
		IDLE 	:	bf0_next_state = ( bf1_current_state == IDLE ) ? WRING : IDLE ;
		WRING 	:	bf0_next_state = (		!write_last		) ? 			WRING	:
										( bf1_current_state == RD_DONE ) ?	READY	: WR_DONE	;
		READY	:	bf0_next_state = RDING ;
		WR_DONE	:	bf0_next_state = ( bf1_current_state==RDING ) ? 		(read_done)? READY : WR_DONE 	: 
										( bf1_current_state==RD_DONE ) ? 	READY : 
											( (bf1_current_state==IDLE) | (bf1_current_state==WRING) ) ? READY : WR_DONE ;
		RDING 	:	bf0_next_state = ( read_done ) ? RD_DONE : RDING ;		//need read last
		RD_DONE :	bf0_next_state = ( bf1_current_state== WRING ) ? RD_DONE : WRING ;

		default: bf0_next_state = IDLE ;
	endcase
end

always @(*) begin
	case (bf1_current_state)
		IDLE 	:	bf1_next_state = ( bf0_current_state == IDLE ) ? IDLE : 
										( (bf0_current_state == WRING) & write_last ) ? WRING : IDLE ;
		WRING 	:	bf1_next_state = (		!write_last		) ? 			WRING	:
										( bf0_current_state == RD_DONE ) ?	READY	: WR_DONE	;
		READY	:	bf1_next_state = RDING ;
		// WR_DONE	:	bf1_next_state = ( read_done ) ? READY : WR_DONE ;
		WR_DONE	:	bf1_next_state = ( bf0_current_state==RDING ) ? 		(read_done)? READY : WR_DONE 	: 
										( bf0_current_state==RD_DONE ) ? 	READY : 
											( (bf0_current_state==IDLE) | (bf0_current_state==WRING) ) ? READY : WR_DONE ;
		RDING 	:	bf1_next_state = ( read_done ) ? RD_DONE : RDING ;		//need read last
		RD_DONE :	bf1_next_state = ( bf0_current_state== WRING ) ? RD_DONE : WRING ;

		default: bf1_next_state = IDLE ;
	endcase
end

// ============================================================================

always @(posedge clk ) begin
	if( reset )begin
		read_start <= 1'd0 ;
	end
	else begin
		if( (bf0_current_state==RDING ) | (bf1_current_state==RDING ))begin
			if( !read_busy )begin
				read_start <= 1'd1 ;
			end
			else begin
				read_start <= 1'd0 ;
			end
		end
		else begin
			read_start <= 1'd0 ;
		end
	end
end

//-----------------------------------------------------------------------------




endmodule