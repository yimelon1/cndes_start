// ============================================================================
// Designer : Yi_Yuan Chen
// Create   : 2022.10.20
// Ver      : 3.0
// Func     : FSM with instruction get testbench, every state need 10 cycle to done
// 			and test for start instruction on different cycle 
// ============================================================================


// `define VIVA
`define End_CYCLE  10000      // Modify cycle times once your design need more cycle times!
`define NI_DELAY  2		// NONIDEAL delay latency

`ifdef RTL
	`timescale 1ns/100ps
    `define CYCLE 5	// 100MHz  1ns*`CYCLE = 10ns / cycle
`endif
`ifdef GATE
	`timescale 1ns/1ps
    `define CYCLE 3.3
`endif
`ifdef VIVA
	`timescale 1ns/100ps
    `define CYCLE 10	// 100MHz
`endif

`ifdef RTL
	`define KER_PAT_0 "../PAT/wsram_pat_0.dat"
	`define KER_PAT_1 "../PAT/wsram_pat_1.dat"
	`define KER_PAT_2 "../PAT/wsram_pat_2.dat"
	`define KER_PAT_3 "../PAT/wsram_pat_3.dat"
	`define KER_PAT_4 "../PAT/wsram_pat_4.dat"
	`define KER_PAT_5 "../PAT/wsram_pat_5.dat"
	`define KER_PAT_6 "../PAT/wsram_pat_6.dat"
	`define KER_PAT_7 "../PAT/wsram_pat_7.dat"
`endif




module fsm_check_tb();
	

	parameter TBITS = 64;
	parameter TBYTE = 8;

	parameter IFMAP_SIZE   = 173056;
	parameter TB_ISRAM_DEPTH	=	300 ;

	localparam IFMAP_SRAM_ADDBITS = 11       ;
	localparam IFMAP_SRAM_DATA_WIDTH = 64    ;
//----------------------------------------------------

//----------------------------------------------------


	reg [30:0] cycle=0;

	reg  clk;         
	reg  reset;       


	logic rstn = 1;
	wire [TBITS-1: 0 ]	isif_data_dout			;
	wire [TBYTE-1: 0 ]	isif_strb_dout			;
	wire 				isif_last_dout			;
	wire 				isif_user_dout			;
	wire 				isif_empty_n			;
	wire 				isif_read				;

	reg              S_AXIS_MM2S_TVALID = 0;
	wire             S_AXIS_MM2S_TREADY;
	reg  [TBITS-1:0] S_AXIS_MM2S_TDATA = 0;
	reg  [TBYTE-1:0] S_AXIS_MM2S_TKEEP = 0;
	reg  [1-1:0]     S_AXIS_MM2S_TLAST = 0;



//---------- pattern declare-----------------
logic tb_memread_done ;
reg    [TBITS-1 : 0]      ifmap        [0:IFMAP_SIZE-1];

logic [63:0] ker_sram_0 [0:2047];
logic [63:0] ker_sram_1 [0:2047];
logic [63:0] ker_sram_2 [0:2047];
logic [63:0] ker_sram_3 [0:2047];
logic [63:0] ker_sram_4 [0:2047];
logic [63:0] ker_sram_5 [0:2047];
logic [63:0] ker_sram_6 [0:2047];
logic [63:0] ker_sram_7 [0:2047];


//--------------------------------------------
//-------------  tb random function test ---------------
	logic [64-1 :0 ] check_ifmaparray0 ;
	logic [64-1 :0 ] check_ifmaparray1 ;
	logic [64-1 :0 ] check_ifmaparray2 ;
	logic [64-1 :0 ] check_ifmaparray3 ;
	logic [64-1 :0 ] check_ifmaparray4 ;
	logic [64-1 :0 ] check_ifmaparray5 ;


integer  iix , i1 , i0 ;



//----------  ker w testbench --------------------
	reg tst_sram_rw;
//----------- test kernel store module ------------------------
	logic ker_write_done;
	logic ker_write_busy;
	logic start_ker_write;
//--------------------------------------------------------------
//----------- test kernel read module ------------------------
	logic ker_read_done;
	logic ker_read_busy;
	logic start_ker_read;
//--------------------------------------------------------------
	logic [63:0] dout_kersr_0 , dout_kersr_1 , dout_kersr_2 , dout_kersr_3 , dout_kersr_4 , dout_kersr_5 , dout_kersr_6 , dout_kersr_7 ;
	logic ksr_valid_0 , ksr_valid_1 , ksr_valid_2 , ksr_valid_3 , ksr_valid_4 , ksr_valid_5 , ksr_valid_6 , ksr_valid_7 ;
	logic ksr_final_0 , ksr_final_1 , ksr_final_2 , ksr_final_3 , ksr_final_4 , ksr_final_5 , ksr_final_6 , ksr_final_7 ;

// testbench data collect
	logic [63:0] dout_kersr_0_dly0 , dout_kersr_1_dly0 , dout_kersr_2_dly0 , dout_kersr_3_dly0 , dout_kersr_4_dly0 , dout_kersr_5_dly0 , dout_kersr_6_dly0 , dout_kersr_7_dly0 ;
	logic ksr_valid_0_dly0 , ksr_valid_1_dly0 , ksr_valid_2_dly0 , ksr_valid_3_dly0 , ksr_valid_4_dly0 , ksr_valid_5_dly0 , ksr_valid_6_dly0 , ksr_valid_7_dly0		;
	logic ksr_final_0_dly0 , ksr_final_1_dly0 , ksr_final_2_dly0 , ksr_final_3_dly0 , ksr_final_4_dly0 , ksr_final_5_dly0 , ksr_final_6_dly0 , ksr_final_7_dly0				;


// =============================================================================
// =======		instance 	===================================================
// =============================================================================

	ker_tset kt001 (
		.clk	(	clk		),
		.reset	(	reset	),

		.ker_write_data_din		(	isif_data_dout	),
		.ker_write_empty_n_din	(	isif_empty_n	),
		.ker_write_read_dout	(	isif_read		),

		.ker_write_done 		(	ker_write_done	),
		.ker_write_busy 		(	ker_write_busy	),
		.start_ker_write		(	start_ker_write	),

		.ker_read_done 			(	ker_read_done 	),
		.ker_read_busy 			(	ker_read_busy 	),
		.start_ker_read			(	start_ker_read	),

		//----generated by ker_top_mod.py------ 
		//----top port list for other module instance------ 
		.dout_kersr_0 ( dout_kersr_0 ), .ksr_valid_0  ( ksr_valid_0 ), .ksr_final_0  ( ksr_final_0 ), //----instance KER top_0---------
		.dout_kersr_1 ( dout_kersr_1 ), .ksr_valid_1  ( ksr_valid_1 ), .ksr_final_1  ( ksr_final_1 ), //----instance KER top_1---------
		.dout_kersr_2 ( dout_kersr_2 ), .ksr_valid_2  ( ksr_valid_2 ), .ksr_final_2  ( ksr_final_2 ), //----instance KER top_2---------
		.dout_kersr_3 ( dout_kersr_3 ), .ksr_valid_3  ( ksr_valid_3 ), .ksr_final_3  ( ksr_final_3 ), //----instance KER top_3---------
		.dout_kersr_4 ( dout_kersr_4 ), .ksr_valid_4  ( ksr_valid_4 ), .ksr_final_4  ( ksr_final_4 ), //----instance KER top_4---------
		.dout_kersr_5 ( dout_kersr_5 ), .ksr_valid_5  ( ksr_valid_5 ), .ksr_final_5  ( ksr_final_5 ), //----instance KER top_5---------
		.dout_kersr_6 ( dout_kersr_6 ), .ksr_valid_6  ( ksr_valid_6 ), .ksr_final_6  ( ksr_final_6 ), //----instance KER top_6---------
		.dout_kersr_7 ( dout_kersr_7 ), .ksr_valid_7  ( ksr_valid_7 ), .ksr_final_7  ( ksr_final_7 ), //----instance KER top_7---------


		.tst_sram_rw			(	tst_sram_rw		)
	
	);

	INPUT_STREAM_if		#(
		.TBITS	(	TBITS	),
		.TBYTE	(	TBYTE	)
	)
	axififo_in (
		// AXI4-Stream singals
		.ACLK       (	clk	),
		.ARESETN    (	rstn	),
		.TVALID     (	S_AXIS_MM2S_TVALID	),
		.TREADY     (	S_AXIS_MM2S_TREADY	),
		.TDATA      (	S_AXIS_MM2S_TDATA	),
		.TKEEP      (	S_AXIS_MM2S_TKEEP	),
		.TLAST      (	S_AXIS_MM2S_TLAST	),
		.TUSER      ( 1'b0 ),

		// User signals
		.isif_data_dout         (	isif_data_dout		),
		.isif_strb_dout         (	isif_strb_dout		),
		.isif_last_dout         (	isif_last_dout		),
		.isif_user_dout         (	isif_user_dout		),
		.isif_empty_n           (	isif_empty_n		),
		.isif_read				(	isif_read			)
	);


// =============================================================================
// ================		random function 		================================
// =============================================================================


	function int unsigned getrand;
		input int unsigned maxvalue ; 
		input int unsigned minvalue ; 
		begin
			getrand = $urandom_range(maxvalue , minvalue);
		end
	endfunction
	//------------- check random ---------------------
	assign check_ifmaparray0	 = getrand(10 , 15) ;
	assign check_ifmaparray1	 = getrand(20 , 50) ;
	assign check_ifmaparray2	 = getrand(20 , 50);
	// assign check_ifmaparray3	 = ifmap[ 180 ] ;
	// assign check_ifmaparray4	 = ifmap[ 240 ] ;
	// assign check_ifmaparray5	 = ifmap[ 560 ] ;
// =============================================================
	


// =============================================================================
// ================		clock generate & end cycle		========================
// =============================================================================

	initial clk = 1;

	always begin #(`CYCLE / 2) clk = ~clk; end
	always@(*)begin
		rstn = ~reset;
	end
	
	always @(posedge clk) begin
		cycle <= cycle+1;
		if (cycle > `End_CYCLE) begin
			$display("********************************************************************");
			$display("**  Failed waiting Valid signal, Simulation STOP at cycle %d **",cycle);
			$display("**  If needed, You can increase End_CYCLE value in tp.v           **");
			$display("********************************************************************");
			$finish;
		end
	end
// =============================================================




// =============================================================================
// ================		fsdb dump +mda+packedmda		========================
// ================		Kernel data load readmemh		========================
// =============================================================================

	initial begin
		`ifdef RTL
			$fsdbDumpfile("tbker.fsdb");
			$fsdbDumpvars(0,"+mda","+packedmda");		//++
			$fsdbDumpMDA();
		`elsif GATE
			$sdf_annotate(`SDFFILE,top_U);
			$fsdbDumpfile("dla_top_SYN.fsdb");
			$fsdbDumpvars();
		`else 
		`endif
	end

	initial begin // initial pattern and expected result
		wait(reset==1);
		tb_memread_done = 0; 
		//--------- pattern reading start -----------
		$readmemh(`KER_PAT_0, ker_sram_0);
		$readmemh(`KER_PAT_1, ker_sram_1);
		$readmemh(`KER_PAT_2, ker_sram_2);
		$readmemh(`KER_PAT_3, ker_sram_3);
		$readmemh(`KER_PAT_4, ker_sram_4);
		$readmemh(`KER_PAT_5, ker_sram_5);
		$readmemh(`KER_PAT_6, ker_sram_6);
		$readmemh(`KER_PAT_7, ker_sram_7);
		//--------- pattern reading end -----------	
		#1;
		tb_memread_done = 1;

	end

// =============================================================



	// -------------- main FSM testing ------------------------

	// -------------- main FSM testing ------------------------

	//start test gi circuit
	initial begin
		#1;
		reset = 0;
		#( `CYCLE*3 ) ;
		reset = 1;
		//-----------reset signal start ------------------
		S_AXIS_MM2S_TKEEP = 'hff;
		S_AXIS_MM2S_TLAST = 0 ;
		start_ker_write = 0;
		start_ker_read = 0 ;
		//-----------reset signal end ------------------
		#( `CYCLE*4 + `NI_DELAY ) ;
		reset = 0;
		#( `CYCLE*5 ) ;


		//----- wait mem read --------------
		wait(tb_memread_done) ;
		#( `CYCLE*5 ) ;
		// //------- ker type1 store start -----------------
		// wait( ker_write_busy==1'd0 );
		// tst_sram_rw = 1 ;
		// @( posedge clk );
		// start_ker_write = 1;
		// #( `CYCLE*3 ) ;
		// @( posedge clk );
		// start_ker_write = 0;

		// for( i0 = 0 ; i0 <8 ; i0 = i0 + 1)begin
		// 	@( posedge clk );
		// 		S_AXIS_MM2S_TLAST = 0 ;
		// 		S_AXIS_MM2S_TVALID = 0 ;
		// 	for( i1=0 ; i1<288 ; i1=i1+1 )begin
		// 		@(posedge clk);
		// 			S_AXIS_MM2S_TVALID=1;
		// 			S_AXIS_MM2S_TDATA = ker_sram_0[ i1  ]	;
		// 			if(  i1==(  287   ) )begin
		// 				S_AXIS_MM2S_TLAST = 1 ;
		// 			end
		// 			wait(S_AXIS_MM2S_TREADY);
		// 	end
		// 	@(posedge clk);
		// 		S_AXIS_MM2S_TVALID = 0 ;
		// 		S_AXIS_MM2S_TLAST = 0 ;
		// 		#(getrand(58 , 15)) ;
		// end
		
		// @(posedge clk);
		// tst_sram_rw = 1 ;
		//------- ker type2 store start -----------------
		wait( ker_write_busy==1'd0 );
		tst_sram_rw = 1 ;
		@( posedge clk );
		start_ker_write = 1;
		#( `CYCLE*3 ) ;
		@( posedge clk );
		start_ker_write = 0;
		
		for( i0 = 0 ; i0 <8 ; i0 = i0 + 1)begin
			@( posedge clk );
				S_AXIS_MM2S_TLAST = 0 ;
				S_AXIS_MM2S_TVALID = 0 ;
			for( i1=0 ; i1<288 ; i1=i1+1 )begin
				@(posedge clk);
					S_AXIS_MM2S_TVALID=1;
					S_AXIS_MM2S_TDATA = ker_sram_0[ i1  ]	;
					if(  (i1==287)    && ( i0 == 7 ) )begin
						S_AXIS_MM2S_TLAST = 1 ;
					end
					wait(S_AXIS_MM2S_TREADY);
			end

		end
		
		@(posedge clk);
			S_AXIS_MM2S_TVALID = 0 ;
			S_AXIS_MM2S_TLAST = 0 ;
			#(getrand(58 , 15)) ;
		@(posedge clk);
		tst_sram_rw = 0 ;

		#(getrand(58 , 15)) ;
		wait( ker_read_busy==1'd0 );
		tst_sram_rw = 0 ;
		@( posedge clk );
		start_ker_read = 1;
		#( `CYCLE*3 ) ;
		@( posedge clk );
		start_ker_read = 0;
		
		#(getrand(58 , 15)) ;
		wait( ker_read_done==1'd1 );




	end 


// =============================================================================
// ================		kernel sram read data check		========================
// =============================================================================
	always @(posedge clk ) begin
		dout_kersr_0_dly0 <= dout_kersr_0 ;
		dout_kersr_1_dly0 <= dout_kersr_1 ;
		dout_kersr_2_dly0 <= dout_kersr_2 ;
		dout_kersr_3_dly0 <= dout_kersr_3 ;
		dout_kersr_4_dly0 <= dout_kersr_4 ;
		dout_kersr_5_dly0 <= dout_kersr_5 ;
		dout_kersr_6_dly0 <= dout_kersr_6 ;
		dout_kersr_7_dly0 <= dout_kersr_7 ;

		ksr_valid_0_dly0 <= ksr_valid_0 ;
		ksr_valid_1_dly0 <= ksr_valid_1 ;
		ksr_valid_2_dly0 <= ksr_valid_2 ;
		ksr_valid_3_dly0 <= ksr_valid_3 ;
		ksr_valid_4_dly0 <= ksr_valid_4 ;
		ksr_valid_5_dly0 <= ksr_valid_5 ;
		ksr_valid_6_dly0 <= ksr_valid_6 ;
		ksr_valid_7_dly0 <= ksr_valid_7 ;

		ksr_final_0_dly0 <= ksr_final_0 ;
		ksr_final_1_dly0 <= ksr_final_1 ;
		ksr_final_2_dly0 <= ksr_final_2 ;
		ksr_final_3_dly0 <= ksr_final_3 ;
		ksr_final_4_dly0 <= ksr_final_4 ;
		ksr_final_5_dly0 <= ksr_final_5 ;
		ksr_final_6_dly0 <= ksr_final_6 ;
		ksr_final_7_dly0 <= ksr_final_7 ;
	end

endmodule