// ============================================================================
// Designer : Yi_Yuan Chen
// Create   : 2022.12.09
// Ver      : 1.0
// Func     : output top module
// ============================================================================
//      Instance Name:              OT_SRAM
//      Words:                      1024
//      Bits:                       64
//      Mux:                        8
//      Drive:                      6
//      Write Mask:                 Off
//      Extra Margin Adjustment:    On
//      Accelerated Retention Test: Off
//      Redundant Rows:             0
//      Redundant Columns:          0
//      Test Muxes                  Off
//----------------------------------------------------------------------------------
//	/----------\     /-----------\     /---------\     /----------\    /---------\
//	| Quan_mod | --> | qtbuf_mod | --> | qtbfifo | --> | ot_write | -->| ot_read |    
//	\----------/     \-----------/     \---------/     \----------/    \---------/
//--------------------------------------------------------------------------------


module ot_top (	
	clk ,
	reset ,

	fifo_full_n		,
	fifo_write		,
	fifo_last		,
	fifo_data		,

	tst_read_last	,
	valid_in 	,
	data_in		


);
	

	localparam SRAM_DATA_BITS = 64;
	localparam SRAM_ADDR_BITS = 10;

//-----------------------------------------------------------------------------

	input clk		;
	input reset		;

	input valid_in 	;
	input [ 8-1 : 0 ]		data_in		;
	input tst_read_last ;

	input 	fifo_full_n		;
	output	fifo_write		;
	output	fifo_last		;
	output [ SRAM_DATA_BITS-1 : 0 ]	fifo_data		;
	
//-----------------------------------------------------------------------------

//----generated by ot_top_mod.py------ 
//---- ot_top declare OT_SRAM start------ 
wire cen_otsr_0 ,cen_otsr_1 ; 
wire wen_otsr_0 ,wen_otsr_1 ; 
wire [ 10 -1 : 0 ] addr_otsr_0 ,addr_otsr_1 ; 
wire [ 64 -1 : 0 ] din_otsr_0 ,din_otsr_1 ; 
wire [ 64 -1 : 0 ] dout_otsr_0 ,dout_otsr_1 ; 
//---- ot top declare OT_SRAM end------ 


//----declare ot_top sram read signal start------ 
wire osr_cen_otsr_0 ; 
wire osr_wen_otsr_0 ; 
wire [ 10 -1 : 0 ] osr_addr_otsr_0 ; 
wire [ 64 -1 : 0 ] osr_dout_otsr_0 ; 
//----declare ot_top sram read signal  end------ 


//----declare ot_top sram write signal start------ 
wire osw_cen_otsr_0 ; 
wire osw_wen_otsr_0 ; 
wire [ 10 -1 : 0 ] osw_addr_otsr_0 ; 
wire [ 64 -1 : 0 ] osw_din_otsr_0 ; 
//----declare ot_top sram write signal  end------ 




localparam BUF_STATE_BITS = 3;
localparam IDLE 	= 3'd0;
localparam READY 	= 3'd1;

localparam WRING 	= 3'd2;
localparam WR_DONE 	= 3'd3;
localparam RDING 	= 3'd4;
localparam RD_DONE 	= 3'd5;

reg [BUF_STATE_BITS-1: 0 ] bf0_current_state ;
reg [BUF_STATE_BITS-1: 0 ] bf0_next_state ;

reg [BUF_STATE_BITS-1: 0 ] bf1_current_state ;
reg [BUF_STATE_BITS-1: 0 ] bf1_next_state ;


wire write_last ;
wire dual_done ;

reg read_start ;
wire read_busy ;
wire read_done ;

//------- qtb and fifo signal --------
wire fifo_empty_n 	;
wire fifo_read 		;
wire valid_to_ot	;
wire [ 64-1 : 0 ]data64_to_ot	;
wire [ 64-1 : 0 ] fifo_data64	;
wire fifo_w_empty_n	;
wire fifo_w_read	;
//-----------------------------------------------------------------------------



// =============================================================================
// ============================		instance		========================
// =============================================================================
//----generated by ot_top_mod.py------ 
//----instance OT_SRAM start------ 
OT_SRAM otbf_0(.Q(	dout_otsr_0 ),	.CLK( clk ),.CEN( cen_otsr_0 ),.WEN( wen_otsr_0 ),.A( addr_otsr_0 ),.D( din_otsr_0 ),.EMA( 3'b0 ));//----instance OT SRAM_0---------
OT_SRAM otbf_1(.Q(	dout_otsr_1 ),	.CLK( clk ),.CEN( cen_otsr_1 ),.WEN( wen_otsr_1 ),.A( addr_otsr_1 ),.D( din_otsr_1 ),.EMA( 3'b0 ));//----instance OT SRAM_1---------
//----instance OT_SRAM end------ 




assign din_otsr_0 	= osw_din_otsr_0 ;
assign cen_otsr_0 	= ( bf0_current_state == WRING )? osw_cen_otsr_0 : 
						( bf0_current_state == RDING )? osr_cen_otsr_0 : 1'd1 	;
assign wen_otsr_0 	= ( bf0_current_state == WRING )? osw_wen_otsr_0 :  1'd1 	;
assign addr_otsr_0	= ( bf0_current_state == WRING )? osw_addr_otsr_0 : 
						( bf0_current_state == RDING )? osr_addr_otsr_0 : 10'd0 	;

assign din_otsr_1 	= osw_din_otsr_0 	;
assign cen_otsr_1 	= ( bf1_current_state == WRING )? osw_cen_otsr_0 : 
						( bf1_current_state == RDING )? osr_cen_otsr_0 : 1'd1 	;
assign wen_otsr_1 	= ( bf1_current_state == WRING )? osw_wen_otsr_0 :  1'd1 	;
assign addr_otsr_1	= ( bf1_current_state == WRING )? osw_addr_otsr_0 : 
						( bf1_current_state == RDING )? osr_addr_otsr_0 : 10'd0 	;


assign osr_dout_otsr_0 = ( bf0_current_state == RDING )? dout_otsr_0 :
							( bf1_current_state == RDING )? dout_otsr_1 :	64'd0 ;




assign fifo_w_empty_n = (  (bf0_current_state == WRING ) | ( bf1_current_state == WRING ) ) ? fifo_empty_n : 1'd0 ;
assign fifo_read = (  (bf0_current_state == WRING ) | ( bf1_current_state == WRING ) ) ? 	fifo_w_read : 1'd0 ;



ot_write #(
	.ADDR_FINAL( 10 )
)ow000 (
	.clk			(	clk				),
	.reset			(	reset			),
	.valid_in 		(	valid_in 		),
	.data_in		(	fifo_data64			),
	.fifo_empty_n	(	fifo_w_empty_n	),
	.fifo_read 		(	fifo_w_read	),

	.last			(	write_last		),
	.cen_otsr		(	osw_cen_otsr_0		),
	.wen_otsr		(	osw_wen_otsr_0		),
	.addr_otsr		(	osw_addr_otsr_0		),
	.data_for_sram	(	osw_din_otsr_0		)

);


ot_read #(
	.ADDR_FINAL( 10 )
)
or111 (
	.clk			(	clk				),
	.reset			(	reset			),

	.start			(	read_start	),
	.busy			(	read_busy	),
	.done			(	read_done	),
	.fifo_full_n	(	fifo_full_n	),
	.fifo_write		(	fifo_write	),
	.fifo_last		(	fifo_last	),
	.fifo_data		(	fifo_data	),

	.data_from_sram	(	osr_dout_otsr_0	),
	.addr_otsr		(	osr_addr_otsr_0	),
	.cen_otsr		(	osr_cen_otsr_0	),
	.wen_otsr		(	osr_wen_otsr_0	)

);


yi_fifo  qtbfifo(
	.clk			(	clk		),
	.reset			(	reset	),
	.valid_in 		(	valid_to_ot	),
	.data_in		(	data64_to_ot	),
	// .error			(		),	// we loss output data cause something wrong
	.empty_n		(	fifo_empty_n	),
	.read			(	fifo_read		),
	.data_out		(	fifo_data64		)
);


ot_qtbuf	qtb00(
	.clk 		(	clk	),
	.reset 		( reset	),
	
	.q_out			(	data_in			),
	.q_valid		(	valid_in		),
	
	.out64bits		(	data64_to_ot	),
	.valid_out		(	valid_to_ot		)

);


// =============================================================================
always @(posedge clk ) begin
	if(reset )begin
		bf0_current_state <= WRING ;
		bf1_current_state <= IDLE ;
	end
	else begin
		bf0_current_state <= bf0_next_state ;
		bf1_current_state <= bf1_next_state ;
	end
end


always @(*) begin
	case (bf0_current_state)
		IDLE 	:	bf0_next_state = ( bf1_current_state == IDLE ) ? WRING : IDLE ;
		WRING 	:	bf0_next_state = (		!write_last		) ? 			WRING	:
										( bf1_current_state == RD_DONE ) ?	READY	: WR_DONE	;
		READY	:	bf0_next_state = RDING ;
		WR_DONE	:	bf0_next_state = ( bf1_current_state==RDING ) ? 		(read_done)? READY : WR_DONE 	: 
										( bf1_current_state==RD_DONE ) ? 	READY : 
											( (bf1_current_state==IDLE) | (bf1_current_state==WRING) ) ? READY : WR_DONE ;
		RDING 	:	bf0_next_state = ( read_done ) ? RD_DONE : RDING ;		//need read last
		RD_DONE :	bf0_next_state = ( bf1_current_state== WRING ) ? RD_DONE : WRING ;

		default: bf0_next_state = IDLE ;
	endcase
end

always @(*) begin
	case (bf1_current_state)
		IDLE 	:	bf1_next_state = ( bf0_current_state == IDLE ) ? IDLE : 
										( (bf0_current_state == WRING) & write_last ) ? WRING : IDLE ;
		WRING 	:	bf1_next_state = (		!write_last		) ? 			WRING	:
										( bf0_current_state == RD_DONE ) ?	READY	: WR_DONE	;
		READY	:	bf1_next_state = RDING ;
		// WR_DONE	:	bf1_next_state = ( read_done ) ? READY : WR_DONE ;
		WR_DONE	:	bf1_next_state = ( bf0_current_state==RDING ) ? 		(read_done)? READY : WR_DONE 	: 
										( bf0_current_state==RD_DONE ) ? 	READY : 
											( (bf0_current_state==IDLE) | (bf0_current_state==WRING) ) ? READY : WR_DONE ;
		RDING 	:	bf1_next_state = ( read_done ) ? RD_DONE : RDING ;		//need read last
		RD_DONE :	bf1_next_state = ( bf0_current_state== WRING ) ? RD_DONE : WRING ;

		default: bf1_next_state = IDLE ;
	endcase
end

// ============================================================================

always @(posedge clk ) begin
	if( reset )begin
		read_start <= 1'd0 ;
	end
	else begin
		if( (bf0_current_state==RDING ) | (bf1_current_state==RDING ))begin
			if( !read_busy )begin
				read_start <= 1'd1 ;
			end
			else begin
				read_start <= 1'd0 ;
			end
		end
		else begin
			read_start <= 1'd0 ;
		end
	end
end


endmodule